`timescale 1 ns/ 1 ns

module alu (src_a, src_b, c, data_out);

input [7:0] src_a, src_b;
input [2:0] c;
output [7:0] data_out;



/* implement here */




endmodule
